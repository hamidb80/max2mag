magic
tech mmi25
timestamp 1692605913
use fet_type_pfet_contacts_all_width_2_0 _0
array 0 7 7560 0 6 7720
timestamp 1108712382
transform 1 0 200 0 1 -430
box -660 -360 900 2360
<< end >>
